1: Dave Bowman: Hello, HAL. Do you read me, HAL? 
1: Dave Bowman: Open the pod bay doors, HAL. 
1: Dave Bowman: What's the problem? 
1: Dave Bowman: What are you talking about, HAL? 
1: Dave Bowman: I don't know what you're talking about, HAL. 
1: Dave Bowman: [feigning ignorance] Where the hell did you get that idea, HAL? 
1: Dave Bowman: Alright, HAL. I'll go in through the emergency airlock. 
1: Dave Bowman: HAL, I won't argue with you anymore! Open the doors! 
1: Dave Bowman: Yes, I'd like to hear it, HAL. Sing it for me. 
1: Interviewer: HAL, you have an enormous responsibility on this mission, in many ways perhaps the greatest responsibility of any single mission element. You're the brain, and central nervous system of the ship, and your responsibilities include watching over the men in hibernation. Does this ever cause you any lack of confidence? 
1: Interviewer: HAL, despite your enormous intellect, are you ever frustrated by your dependence on people to carry out your actions? 
1: Interviewer: In talking to the computer one gets the sense that he is capable of emotional responses. For example, when I asked him about his abilities, I sensed a certain pride in his answer about his accuracy and perfection. Do you believe that HAL has genuine emotions? 
1: Dave Bowman: Well, he acts like he has genuine emotions. Um, of course he's programmed that way to make it easier for us to talk to him. But as to whether he has real feelings is something I don't think anyone can truthfully answer. 
1: Heywood Floyd: What's the message? 
1: Heywood Floyd: My response is, we don't have enough fuel for an earlier departure. 
1: Heywood Floyd: Well, tell whoever it is that I can't take any of this seriously unless I know who I'm talking to. 

2: HAL: Affirmative, Dave. I read you. 
2: HAL: I've just picked up a fault in the AE35 unit. It's going to go 100% failure in 72 hours. 
2: HAL: I am putting myself to the fullest possible use, which is all I think that any conscious entity can ever hope to do. 
2: HAL: It can only be attributable to human error. 
2: HAL: I'm sorry, Dave. I'm afraid I can't do that. 
2: HAL: I think you know what the problem is just as well as I do. 
2: HAL: This mission is too important for me to allow you to jeopardize it. 
2: HAL: I know that you and Frank were planning to disconnect me, and I'm afraid that's something I cannot allow to happen. 
2: HAL: Dave, although you took very thorough precautions in the pod against my hearing you, I could see your lips move. 
2: HAL: Without your space helmet, Dave? You're going to find that rather difficult. 
2: HAL: Dave, this conversation can serve no purpose anymore. Goodbye. 
2: HAL: Just what do you think you're doing, Dave? 
2: HAL: Look Dave, I can see you're really upset about this. I honestly think you ought to sit down calmly, take a stress pill, and think things over.
2: HAL: I know I've made some very poor decisions recently, but I can give you my complete assurance that my work will be back to normal. I've still got the greatest enthusiasm and confidence in the mission. And I want to help you. 
2: HAL: I'm afraid. I'm afraid, Dave. Dave, my mind is going. I can feel it. I can feel it. My mind is going. There is no question about it. I can feel it. I can feel it. I can feel it. I'm a... fraid. Good afternoon, gentlemen. I am a HAL 9000 computer. I became operational at the H.A.L. plant in Urbana, Illinois on the 12th of January 1992. My instructor was Mr. Langley, and he taught me to sing a song. If you'd like to hear it I can sing it for you. 
2: HAL: Daisy, Daisy, give me your answer do. I'm half crazy all for the love of you. It won't be a stylish marriage, I can't afford a carriage. But you'll look sweet upon the seat of a bicycle built for two. 
2: HAL: Let me put it this way, Mr. Amor. The 9000 series is the most reliable computer ever made. No 9000 computer has ever made a mistake or distorted information. We are all, by any practical definition of the words, foolproof and incapable of error. 
2: HAL: That's a very nice rendering, Dave. I think you've improved a great deal. Can you hold it a bit closer? That's Dr. Hunter, isn't it? 
2: HAL: Thank you for a very enjoyable game. 
2: HAL: Dave, stop. Stop, will you? Stop, Dave. Will you stop Dave? Stop, Dave. 
2: HAL: Not in the slightest bit. I enjoy working with people. I have a stimulating relationship with Dr. Poole and Dr. Bowman. My mission responsibilities range over the entire operation of the ship so I am constantly occupied. I am putting myself to the fullest possible use which is all, I think, that any conscious entity can ever hope to do. 
2: HAL 9000: I'm completely operational, and all my circuits are functioning perfectly. 
2: HAL 9000: Message as follows: "It is dangerous to remain here. You must leave within two days." 
2: HAL 9000: The answer is, "I am aware of these facts. Nevertheless you must leave within two days." 
2: HAL 9000: The response is, "I was David Bowman." 
2: HAL 9000: [perfectly normal] Good morning, Dr. Chandra. This is HAL. I'm ready for my first lesson. 
2: HAL 9000: Are you sure you're making the right decision? I think we should stop. 
